`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07/04/2024 09:12:52 AM
// Design Name: 
// Module Name: sbox5
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module sbox5(
       input logic [5:0] X,
       output logic [3:0] Y
    );
    
     assign Y =  (X == 6'b0_0000_0) ? 4'd2 :
                (X == 6'b0_0001_0) ? 4'd12 :
                (X==6'b0_0010_0) ? 4'd4 :
                (X==6'b0_0011_0) ? 4'd1 :
                (X==6'b0_0100_0) ? 4'd7 :
                (X==6'b0_0101_0) ? 4'd10 :
                (X==6'b0_0110_0) ? 4'd11 :
                (X==6'b0_0111_0) ? 4'd6 :
                (X==6'b0_1000_0) ? 4'd8  :
                (X==6'b0_1001_0) ? 4'd5 :
                (X==6'b0_1010_0) ? 4'd3  :
                (X==6'b0_1011_0) ? 4'd15 :
                (X==6'b0_1100_0) ? 4'd13 :
                (X==6'b0_1101_0) ? 4'd0 :
                (X==6'b0_1110_0) ? 4'd14 :
                (X==6'b0_1111_0) ? 4'd9 :

                (X == 6'b0_0000_1) ? 4'd14 :
                (X == 6'b0_0001_1) ? 4'd11 :
                (X==6'b0_0010_1) ? 4'd2  :
                (X==6'b0_0011_1) ? 4'd12 :
                (X==6'b0_0100_1) ? 4'd4 :
                (X==6'b0_0101_1) ? 4'd7 :
                (X==6'b0_0110_1) ? 4'd13 :
                (X==6'b0_0111_1) ? 4'd1 :
                (X==6'b0_1000_1) ? 4'd5 :
                (X==6'b0_1001_1) ? 4'd0 :
                (X==6'b0_1010_1) ? 4'd15  :
                (X==6'b0_1011_1) ? 4'd10 :
                (X==6'b0_1100_1) ? 4'd3 :
                (X==6'b0_1101_1) ? 4'd9 :
                (X==6'b0_1110_1) ? 4'd8 :
                (X==6'b0_1111_1) ? 4'd6 :

                (X == 6'b1_0000_0) ? 4'd4 :
                (X == 6'b1_0001_0) ? 4'd2  :
                (X==6'b1_0010_0) ? 4'd1 :
                (X==6'b1_0011_0) ? 4'd11 :
                (X==6'b1_0100_0) ? 4'd10 :
                (X==6'b1_0101_0) ? 4'd13 :
                (X==6'b1_0110_0) ? 4'd7 :
                (X==6'b1_0111_0) ? 4'd8 :
                (X==6'b1_1000_0) ? 4'd15 :
                (X==6'b1_1001_0) ? 4'd9 :
                (X==6'b1_1010_0) ? 4'd12  :
                (X==6'b1_1011_0) ? 4'd5 :
                (X==6'b1_1100_0) ? 4'd6 :
                (X==6'b1_1101_0) ? 4'd3 :
                (X==6'b1_1110_0) ? 4'd0 :
                (X==6'b1_1111_0) ? 4'd14 :

                (X == 6'b1_0000_1) ? 4'd11 :
                (X == 6'b1_0001_1) ? 4'd8 :
                (X==6'b1_0010_1) ? 4'd12 :
                (X==6'b1_0011_1) ? 4'd7 :
                (X==6'b1_0100_1) ? 4'd1 :
                (X==6'b1_0101_1) ? 4'd14 :
                (X==6'b1_0110_1) ? 4'd2 :
                (X==6'b1_0111_1) ? 4'd13 :
                (X==6'b1_1000_1) ? 4'd6 :
                (X==6'b1_1001_1) ? 4'd15 :
                (X==6'b1_1010_1) ? 4'd0 :
                (X==6'b1_1011_1) ? 4'd9 :
                (X==6'b1_1100_1) ? 4'd10 :
                (X==6'b1_1101_1) ? 4'd4 :
                (X==6'b1_1110_1) ? 4'd5 :
                (X==6'b1_1111_1) ? 4'd3 :

                                   4'dX ;


endmodule
